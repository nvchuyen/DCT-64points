module test_DCT1D8P();

reg clk;
reg [3:0] cnt_clk;
reg [23:0] a0, a1, a2, a3, a4, a5, a6, a7;
wire [23:0] w0, w1, w2, w3, w4, w5, w6, w7;
localparam CNT_Clk = 1;

DCT1D8P #(.CNT_Clk(CNT_Clk)) P (.clk(clk),.clk_cnt(cnt_clk),.a0(a0),.a1(a1),.a2(a2),.a3(a3),.a4(a4),.a5(a5),.a6(a6),.a7(a7),
.o0(w0),.o1(w1),.o2(w2),.o3(w3),.o4(w4),.o5(w5),.o6(w6),.o7(w7));

initial
begin
 clk = 1;
 forever  #5 clk = ~clk;
end

initial
begin 
	a0 =  24'b00010111011100101101;//24'b00001000001000000000;
	a1 = 	24'b00010111110110001111;//24'b00001000010000000000;
	a2 =  24'b00011000001010000110;//24'b00001000010000000000;
	a3 =  24'b00011000000111010001;//24'b00001000000100000000;
	a4 =  24'b00011000011100100010;//24'b00001000010100000000;
	a5 =  24'b00011000000011000000;//24'b00001000010100000000;
	a6 =  24'b00011000011000010010;//24'b00001000011000000000;
	a7 =  24'b00011000011111011000;//24'b00001000011100000000;
	#10;
	cnt_clk = 1;
	#10;
	cnt_clk = 2;
	#10;
	cnt_clk = 3;
end 
endmodule  
