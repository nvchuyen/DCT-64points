module testB_DCT1D();

	reg	 clk;
	reg [3:0] cnt_clk;
	reg [23:0] a0,a1,a2,a3,a4,a5,a6,a7;
	reg [23:0] a8,a9,a10,a11,a12,a13,a14,a15;
	reg [23:0] a16,a17,a18,a19,a20,a21,a22,a23;
	reg [23:0] a24,a25,a26,a27,a28,a29,a30,a31;
	reg [23:0] a32,a33,a34,a35,a36,a37,a38,a39;
	reg [23:0] a40,a41,a42,a43,a44,a45,a46,a47;
	reg [23:0] a48,a49,a50,a51,a52,a53,a54,a55;
	reg [23:0] a56,a57,a58,a59,a60,a61,a62,a63;
	wire [23:0] w0,w1,w2,w3,w4,w5,w6,w7;
	wire [23:0] w8,w9,w10,w11,w12,w13,w14,w15;
	wire [23:0] w16,w17,w18,w19,w20,w21,w22,w23;
	wire [23:0] w24,w25,w26,w27,w28,w29,w30,w31;
	wire [23:0] w32,w33,w34,w35,w36,w37,w38,w39;
	wire [23:0] w40,w41,w42,w43,w44,w45,w46,w47;
	wire [23:0] w48,w49,w50,w51,w52,w53,w54,w55;
	wire [23:0] w56,w57,w58,w59,w60,w61,w62,w63;
	localparam CNT_Clk= 1;
	
DCT1D #(.CNT_CLK(CNT_Clk)) testB_DCT2D (.clk(clk),.clk_cnt(cnt_clk),
.a0(a0),.a1(a1),.a2(a2),.a3(a3),.a4(a4),.a5(a5),.a6(a6),.a7(a7),
.a8(a8),.a9(a9),.a10(a10),.a11(a11),.a12(a12),.a13(a13),.a14(a14),.a15(a15),
.a16(a16),.a17(a17),.a18(a18),.a19(a19),.a20(a20),.a21(a21),.a22(a22),.a23(a23),
.a24(a24),.a25(a25),.a26(a26),.a27(a27),.a28(a28),.a29(a29),.a30(a30),.a31(a31),
.a32(a32),.a33(a33),.a34(a34),.a35(a35),.a36(a36),.a37(a37),.a38(a38),.a39(a39),
.a40(a40),.a41(a41),.a42(a42),.a43(a43),.a44(a44),.a45(a45),.a46(a46),.a47(a47),
.a48(a48),.a49(a49),.a50(a50),.a51(a51),.a52(a52),.a53(a53),.a54(a54),.a55(a55),
.a56(a56),.a57(a57),.a58(a58),.a59(a59),.a60(a60),.a61(a61),.a62(a62),.a63(a63),
.o0(w0),.o1(w1),.o2(w2),.o3(w3),.o4(w4),.o5(w5),.o6(w6),.o7(w7),
.o8(w8),.o9(w9),.o10(w10),.o11(w11),.o12(w12),.o13(w13),.o14(w14),.o15(w15),
.o16(w16),.o17(w17),.o18(w18),.o19(w19),.o20(w20),.o21(w21),.o22(w22),.o23(w23),
.o24(w24),.o25(w25),.o26(w26),.o27(w27),.o28(w28),.o29(w29),.o30(w30),.o31(w31),
.o32(w32),.o33(w33),.o34(w34),.o35(w35),.o36(w36),.o37(w37),.o38(w38),.o39(w39),
.o40(w40),.o41(w41),.o42(w42),.o43(w43),.o44(w44),.o45(w45),.o46(w46),.o47(w47),
.o48(w48),.o49(w49),.o50(w50),.o51(w51),.o52(w52),.o53(w53),.o54(w54),.o55(w55),
.o56(w56),.o57(w57),.o58(w58),.o59(w59),.o60(w60),.o61(w61),.o62(w62),.o63(w63));					
	
initial 
begin
	clk =0;
	forever #5 clk = ~clk;
end 

initial 
begin
	a0 = 24'b1000001000000000;//130
	a1 = 24'b1000010000000000;
	a2 = 24'b1000010000000000;
	a3 =  24'b1000000100000000;
	a4 =  24'b1000010100000000;
	a5 =  24'b1000010100000000;
	a6 =  24'b1000011000000000;
	a7 =  24'b1000011100000000;
	
	a8 =  24'b1000011100000000;
	a9 =  24'b1000010100000000;
	a10  =  24'b1000010100000000;
	a11  =  24'b1000001100000000;
	a12 =  24'b1000010100000000;
	a13 =  24'b1000100100000000;
	a14 =  24'b1000101000000000;
	a15 =  24'b1000100000000000;
	
	a16 =  24'b1000010000000000;
	a17 =  24'b1000011000000000;
	a18 =  24'b1000010100000000;
	a19 =  24'b1000100000000000;
	a20 =  24'b1000101100000000;
	a21 =  24'b1000111000000000;
	a22 =  24'b1000100100000000;
	a23 =  24'b1000100100000000;
	
	a24 =  24'b1000100100000000;
	a25 =  24'b1000100000000000;
	a26 =  24'b1000100000000000;
	a27 =  24'b1000011100000000;
	a28 =  24'b1000011100000000;
	a29 =  24'b1000100000000000;
	a30 =  24'b1000011100000000;
	a31 =  24'b1000101000000000;
	
	a32 =  24'b1000101100000000;
	a33 =  24'b1000101000000000;
	a34 =  24'b1000101100000000;
	a35 =  24'b1000011100000000;
	a36 =  24'b1000100000000000;
	a37 =  24'b1000101100000000;
	a38 =  24'b1000100100000000;
	a39 =  24'b1000110000000000;
	
	a40 =  24'b1000011000000000;
	a41 =  24'b1000100000000000;
	a42 =  24'b1000100100000000;
	a43 =  24'b1000100000000000;
	a44 =  24'b1000011000000000;
	a45 =  24'b1000100000000000;
	a46 =  24'b1000100000000000;
	a47 =  24'b1000100000000000;
	
	a48 =  24'b1000100000000000;
	a49 =  24'b1000010100000000;
	a50 =  24'b1000101000000000;
	a51 =  24'b1000100000000000;
	a52 =  24'b1000100000000000;
	a53 =  24'b1000100000000000;
	a54 =  24'b1000101100000000;
	a55 =  24'b1001001000000000;

	
	a56 =  24'b1000101100000000;
	a57 =  24'b1000100100000000;
	a58 =  24'b1000101000000000;
	a59 =  24'b1000011000000000;
	a60 =  24'b1000010100000000;
	a61 =  24'b1000101000000000;
	a62 =  24'b1000110000000000;
	a63 =  24'b1001001000000000;
	
	#10;
	cnt_clk = 1;
	#10;
	cnt_clk = 2;
	#10;
	cnt_clk = 3;
	#10;
	cnt_clk = 4;
	#10;
	cnt_clk = 5;
end 
endmodule 