module DCT2D
(
	input clk, reset,
	input [23:0] a0,a1,a2,a3,a4,a5,a6,a7,
	input [23:0] a8,a9,a10,a11,a12,a13,a14,a15,
	input [23:0] a16,a17,a18,a19,a20,a21,a22,a23,
	input [23:0] a24,a25,a26,a27,a28,a29,a30,a31,
	input [23:0] a32,a33,a34,a35,a36,a37,a38,a39,
	input [23:0] a40,a41,a42,a43,a44,a45,a46,a47,
	input [23:0] a48,a49,a50,a51,a52,a53,a54,a55,
	input [23:0] a56,a57,a58,a59,a60,a61,a62,a63,
	output wire [23:0] o0,o1,o2,o3,o4,o5,o6,o7,
	output wire [23:0] o8,o9,o10,o11,o12,o13,o14,o15,
	output wire [23:0] o16,o17,o18,o19,o20,o21,o22,o23,
	output wire [23:0] o24,o25,o26,o27,o28,o29,o30,o31,
	output wire [23:0] o32,o33,o34,o35,o36,o37,o38,o39,
	output wire [23:0] o40,o41,o42,o43,o44,o45,o46,o47,
	output wire [23:0] o48,o49,o50,o51,o52,o53,o54,o55,
	output wire [23:0] o56,o57,o58,o59,o60,o61,o62,o63
);
localparam size_cnt = 3;
localparam clk_DD1 = 1, clk_DD2 = 5; 
wire [23:0] w0,w1,w2,w3,w4,w5,w6,w7;
wire [23:0] w8,w9,w10,w11,w12,w13,w14,w15;
wire [23:0] w16,w17,w18,w19,w20,w21,w22,w23;
wire [23:0] w24,w25,w26,w27,w28,w29,w30,w31;
wire [23:0] w32,w33,w34,w35,w36,w37,w38,w39;
wire [23:0] w40,w41,w42,w43,w44,w45,w46,w47;
wire [23:0] w48,w49,w50,w51,w52,w53,w54,w55;
wire [23:0] w56,w57,w58,w59,w60,w61,w62,w63;
wire [3:0] cnt_clk;

Cnt_clk 	#(.SIZE_CNT(size_cnt))   cnt_clk1 	(.clk(clk),.reset(reset),.Cnt(cnt_clk));

DCT1D #(.CNT_CLK(clk_DD1)) DD1 (.clk(clk),.clk_cnt(cnt_clk),
.a0(a0),.a1(a1),.a2(a2),.a3(a3),.a4(a4),.a5(a5),.a6(a6),.a7(a7),
.a8(a8),.a9(a9),.a10(a10),.a11(a11),.a12(a12),.a13(a13),.a14(a14),.a15(a15),
.a16(a16),.a17(a17),.a18(a18),.a19(a19),.a20(a20),.a21(a21),.a22(a22),.a23(a23),
.a24(a24),.a25(a25),.a26(a26),.a27(a27),.a28(a28),.a29(a29),.a30(a30),.a31(a31),
.a32(a32),.a33(a33),.a34(a34),.a35(a35),.a36(a36),.a37(a37),.a38(a38),.a39(a39),
.a40(a40),.a41(a41),.a42(a42),.a43(a43),.a44(a44),.a45(a45),.a46(a46),.a47(a47),
.a48(a48),.a49(a49),.a50(a50),.a51(a51),.a52(a52),.a53(a53),.a54(a54),.a55(a55),
.a56(a56),.a57(a57),.a58(a58),.a59(a59),.a60(a60),.a61(a61),.a62(a62),.a63(a63),
.o0(w0),.o1(w1),.o2(w2),.o3(w3),.o4(w4),.o5(w5),.o6(w6),.o7(w7),
.o8(w8),.o9(w9),.o10(w10),.o11(w11),.o12(w12),.o13(w13),.o14(w14),.o15(w15),
.o16(w16),.o17(w17),.o18(w18),.o19(w19),.o20(w20),.o21(w21),.o22(w22),.o23(w23),
.o24(w24),.o25(w25),.o26(w26),.o27(w27),.o28(w28),.o29(w29),.o30(w30),.o31(w31),
.o32(w32),.o33(w33),.o34(w34),.o35(w35),.o36(w36),.o37(w37),.o38(w38),.o39(w39),
.o40(w40),.o41(w41),.o42(w42),.o43(w43),.o44(w44),.o45(w45),.o46(w46),.o47(w47),
.o48(w48),.o49(w49),.o50(w50),.o51(w51),.o52(w52),.o53(w53),.o54(w54),.o55(w55),
.o56(w56),.o57(w57),.o58(w58),.o59(w59),.o60(w60),.o61(w61),.o62(w62),.o63(w63));

DCT1D #(.CNT_CLK(clk_DD2)) DD2 (.clk(clk),.clk_cnt(cnt_clk),
.a0(w0),.a1(w1),.a2(w2),.a3(w3),.a4(w4),.a5(w5),.a6(w6),.a7(w7),
.a8(w8),.a9(w9),.a10(w10),.a11(w11),.a12(w12),.a13(w13),.a14(w14),.a15(w15),
.a16(w16),.a17(w17),.a18(w18),.a19(w19),.a20(w20),.a21(w21),.a22(w22),.a23(w23),
.a24(w24),.a25(w25),.a26(w26),.a27(w27),.a28(w28),.a29(w29),.a30(w30),.a31(w31),
.a32(w32),.a33(w33),.a34(w34),.a35(w35),.a36(w36),.a37(w37),.a38(w38),.a39(w39),
.a40(w40),.a41(w41),.a42(w42),.a43(w43),.a44(w44),.a45(w45),.a46(w46),.a47(w47),
.a48(w48),.a49(w49),.a50(w50),.a51(w51),.a52(w52),.a53(w53),.a54(w54),.a55(w55),
.a56(w56),.a57(w57),.a58(w58),.a59(w59),.a60(w60),.a61(w61),.a62(w62),.a63(w63),
.o0(o0),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.o5(o5),.o6(o6),.o7(o7),
.o8(o8),.o9(o9),.o10(o10),.o11(o11),.o12(o12),.o13(o13),.o14(o14),.o15(o15),
.o16(o16),.o17(o17),.o18(o18),.o19(o19),.o20(o20),.o21(o21),.o22(o22),.o23(o23),
.o24(o24),.o25(o25),.o26(o26),.o27(o27),.o28(o28),.o29(o29),.o30(o30),.o31(o31),
.o32(o32),.o33(o33),.o34(o34),.o35(o35),.o36(o36),.o37(o37),.o38(o38),.o39(o39),
.o40(o40),.o41(o41),.o42(o42),.o43(o43),.o44(o44),.o45(o45),.o46(o46),.o47(o47),
.o48(o48),.o49(o49),.o50(o50),.o51(o51),.o52(o52),.o53(o53),.o54(o54),.o55(o55),
.o56(o56),.o57(o57),.o58(o58),.o59(o59),.o60(o60),.o61(o61),.o62(o62),.o63(o63)
);

endmodule 



